//VIRTUAL_SEQUENCE

