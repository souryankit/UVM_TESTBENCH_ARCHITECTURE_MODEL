//VIRTUAL_SEQUENCER

